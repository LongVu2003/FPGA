`timescale 1ns/1ps
module TB_Mul4x4_4x2matrix;
	reg signed [15:0] A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15;
	reg signed [15:0] B0,B1,B2,B3,B4,B5,B6,B7;
	wire signed [15:0] S0,S1,S2,S3,S4,S5,S6,S7;
	
	Mul4x4_4x2matrix m1(A0,A1,A2,A3,A4,A5,A6,A7,A8,A9,A10,A11,A12,A13,A14,A15,
							B0,B1,B2,B3,B4,B5,B6,B7,
							S0,S1,S2,S3,S4,S5,S6,S7);	
							
	initial begin
		//_____________INIT___________________
		A0  <= 0; A1  <= 0; A2  <= 0; A3  <= 0;
		A4  <= 0; A5  <= 0; A6  <= 0; A7  <= 0;
		A8  <= 0; A9  <= 0; A10 <= 0; A11 <= 0;
		A12 <= 0; A13 <= 0; A14 <= 0; A15 <= 0;
		B1  <= 0; B3  <= 0; B5  <= 0; B7  <= 0;
		B0  <= 0; B2  <= 0; B4  <= 0; B6  <= 0;
		#5
		//_____________TEST1___________________
		/*
			 0.5	 1.5	-1.5	-1.5				-3.5	-3.5
			 0.5	-3.5	-1.5	-1.5    x    	-3.5	-3.5  
			-1.5	 1.5	-3.5	 1.5				 0.5	-3.5
			-3.5	-3.5	 0.5	-3.5				-3.5	-3.5

		*/
		A0  <= 16'h0080; A1  <= 16'h0180; A2  <= 16'hfe80; A3  <= 16'hfe80;
		A4  <= 16'h0080; A5  <= 16'hfc80; A6  <= 16'hfe80; A7  <= 16'hfe80;
		A8  <= 16'hfe80; A9  <= 16'h0180; A10 <= 16'hfc80; A11 <= 16'h0180;
		A12 <= 16'hfc80; A13 <= 16'hfc80; A14 <= 16'h0080; A15 <= 16'hfc80;
		B1  <= 16'hfc80; B3  <= 16'hfc80; B5  <= 16'hfc80; B7  <= 16'hfc80;
		B0  <= 16'hfc80; B2  <= 16'hfc80; B4  <= 16'h0080; B6  <= 16'hfc80;
		
		#5 display;
		
		//_____________TEST2___________________
		/*
			 0.5	 1.5	-1.5	-1.5				-1	 -1
			 0.5	-3.5	-1.5	-1.5    x    	 1	 -2  
			-1.5	 1.5	-3.5	 1.5				 1	 -1
			-3.5	-3.5	 0.5	-3.5				 1	 -1

		*/
		A0  <= 16'h0080; A1  <= 16'h0180; A2  <= 16'hfe80; A3  <= 16'hfe80;
		A4  <= 16'h0080; A5  <= 16'hfc80; A6  <= 16'hfe80; A7  <= 16'hfe80;
		A8  <= 16'hfe80; A9  <= 16'h0180; A10 <= 16'hfc80; A11 <= 16'h0180;
		A12 <= 16'hfc80; A13 <= 16'hfc80; A14 <= 16'h0080; A15 <= 16'hfc80;
		B1  <= 16'hff00; B3  <= 16'hfe00; B5  <= 16'hff00; B7  <= 16'hff00;
		B0  <= 16'hff00; B2  <= 16'h0100; B4  <= 16'h0100; B6  <= 16'h0100;
		
		#5 display;
		
		
		//_____________TEST3___________________
		/*
			 0.5	 1.5	-1.5	-1.5				-1	 -1
			 0.5	-3.5	-1.5	-1.5    x    	 1	 -2  
			-1.5	 1.5	-3.5	 1.5				 1	 -1
			-3.5	-3.5	 0.5	-3.5				 3	 -1

		*/
		A0  <= 16'h0080; A1  <= 16'h0180; A2  <= 16'hfe80; A3  <= 16'hfe80;
		A4  <= 16'h0080; A5  <= 16'hfc80; A6  <= 16'hfe80; A7  <= 16'hfe80;
		A8  <= 16'hfe80; A9  <= 16'h0180; A10 <= 16'hfc80; A11 <= 16'h0180;
		A12 <= 16'hfc80; A13 <= 16'hfc80; A14 <= 16'h0080; A15 <= 16'hfc80;
		B1  <= 16'hff00; B3  <= 16'hfe00; B5  <= 16'hff00; B7  <= 16'hff00;
		B0  <= 16'hff00; B2  <= 16'h0100; B4  <= 16'h0100; B6  <= 16'h0300;
		
		#5 display;
		

		
		
		end
		
		
		task display;
			begin
				$display("Ma tran A");
				$display("[%h %h %h %h]", A0,A1,A2,A3);
				$display("[%h %h %h %h]", A4,A5,A6,A7);
				$display("[%h %h %h %h]", A8,A9,A10,A11);
				$display("[%h %h %h %h]", A12,A13,A14,A15);
				$display("Ma tran B ");
				$display("[%h %h]", B0,B1);
				$display("[%h %h]", B2,B3);
				$display("[%h %h]", B4,B5);
				$display("[%h %h]", B6,B7);
				$display("Ma tran ket qua");
				$display("[%h %h]", S0,S1);
				$display("[%h %h]", S2,S3);
				$display("[%h %h]", S4,S5);
				$display("[%h %h]", S6,S7);
			end
		endtask
endmodule
					
		